<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-61.8331,-330.708,233.765,-476.816</PageViewport>
<gate>
<ID>194</ID>
<type>AE_DFF_LOW</type>
<position>28,-387</position>
<input>
<ID>IN_0</ID>108 </input>
<output>
<ID>OUTINV_0</ID>104 </output>
<output>
<ID>OUT_0</ID>103 </output>
<input>
<ID>clock</ID>105 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2</ID>
<type>AA_LABEL</type>
<position>13,6</position>
<gparam>LABEL_TEXT SR latch using nand gate</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>196</ID>
<type>GA_LED</type>
<position>36,-385</position>
<input>
<ID>N_in0</ID>103 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>197</ID>
<type>GA_LED</type>
<position>36,-388</position>
<input>
<ID>N_in0</ID>104 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>-10.5,-5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>198</ID>
<type>BB_CLOCK</type>
<position>17.5,-391</position>
<output>
<ID>CLK</ID>105 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>5</ID>
<type>AA_TOGGLE</type>
<position>-10.5,-15.5</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>200</ID>
<type>AA_AND2</type>
<position>1.5,-384</position>
<input>
<ID>IN_0</ID>103 </input>
<input>
<ID>IN_1</ID>109 </input>
<output>
<ID>OUT</ID>106 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7</ID>
<type>GA_LED</type>
<position>30.5,-6</position>
<input>
<ID>N_in0</ID>6 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>201</ID>
<type>AA_AND2</type>
<position>1.5,-391.5</position>
<input>
<ID>IN_0</ID>110 </input>
<input>
<ID>IN_1</ID>104 </input>
<output>
<ID>OUT</ID>107 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8</ID>
<type>GA_LED</type>
<position>30,-14.5</position>
<input>
<ID>N_in0</ID>7 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>203</ID>
<type>AE_OR2</type>
<position>10,-387</position>
<input>
<ID>IN_0</ID>106 </input>
<input>
<ID>IN_1</ID>107 </input>
<output>
<ID>OUT</ID>108 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>10</ID>
<type>BA_NAND2</type>
<position>1.5,-6</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>7 </input>
<output>
<ID>OUT</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>11</ID>
<type>BA_NAND2</type>
<position>1.5,-14.5</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>5 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>205</ID>
<type>AA_TOGGLE</type>
<position>-7.5,-385</position>
<output>
<ID>OUT_0</ID>109 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>206</ID>
<type>AA_TOGGLE</type>
<position>-7.5,-390.5</position>
<output>
<ID>OUT_0</ID>110 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>207</ID>
<type>AA_LABEL</type>
<position>-11,-390</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>208</ID>
<type>AA_LABEL</type>
<position>-11,-384.5</position>
<gparam>LABEL_TEXT R</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>209</ID>
<type>AE_DFF_LOW</type>
<position>28,-415.5</position>
<input>
<ID>IN_0</ID>116 </input>
<output>
<ID>OUTINV_0</ID>112 </output>
<output>
<ID>OUT_0</ID>111 </output>
<input>
<ID>clock</ID>113 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_LABEL</type>
<position>37.5,-5.5</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>210</ID>
<type>GA_LED</type>
<position>36,-413.5</position>
<input>
<ID>N_in0</ID>111 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>17</ID>
<type>AA_LABEL</type>
<position>38.5,-14.5</position>
<gparam>LABEL_TEXT Q'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>211</ID>
<type>GA_LED</type>
<position>36,-416.5</position>
<input>
<ID>N_in0</ID>112 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>18</ID>
<type>AA_LABEL</type>
<position>13,-28</position>
<gparam>LABEL_TEXT SR latch using NOR gate</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>212</ID>
<type>BB_CLOCK</type>
<position>17.5,-419.5</position>
<output>
<ID>CLK</ID>113 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>19</ID>
<type>AA_LABEL</type>
<position>-14.5,-4.5</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>213</ID>
<type>AA_AND2</type>
<position>1.5,-412.5</position>
<input>
<ID>IN_0</ID>111 </input>
<input>
<ID>IN_1</ID>117 </input>
<output>
<ID>OUT</ID>114 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_LABEL</type>
<position>-14.5,-15</position>
<gparam>LABEL_TEXT R</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>214</ID>
<type>AA_AND2</type>
<position>1.5,-420</position>
<input>
<ID>IN_0</ID>118 </input>
<input>
<ID>IN_1</ID>112 </input>
<output>
<ID>OUT</ID>115 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>21</ID>
<type>AA_TOGGLE</type>
<position>-8,-39</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>215</ID>
<type>AE_OR2</type>
<position>10,-415.5</position>
<input>
<ID>IN_0</ID>114 </input>
<input>
<ID>IN_1</ID>115 </input>
<output>
<ID>OUT</ID>116 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_TOGGLE</type>
<position>-8,-49.5</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>216</ID>
<type>AA_TOGGLE</type>
<position>-7.5,-413.5</position>
<output>
<ID>OUT_0</ID>117 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>23</ID>
<type>AA_LABEL</type>
<position>-12,-38.5</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>217</ID>
<type>AA_TOGGLE</type>
<position>-7.5,-419</position>
<output>
<ID>OUT_0</ID>118 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_LABEL</type>
<position>-12,-49</position>
<gparam>LABEL_TEXT R</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>218</ID>
<type>AA_LABEL</type>
<position>-11,-418.5</position>
<gparam>LABEL_TEXT J</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>25</ID>
<type>GA_LED</type>
<position>32.5,-40</position>
<input>
<ID>N_in0</ID>11 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>219</ID>
<type>AA_LABEL</type>
<position>-11,-413</position>
<gparam>LABEL_TEXT K</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>26</ID>
<type>GA_LED</type>
<position>32.5,-48.5</position>
<input>
<ID>N_in0</ID>10 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>220</ID>
<type>AA_LABEL</type>
<position>7.5,-401</position>
<gparam>LABEL_TEXT T to JK  Flip Flop</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>27</ID>
<type>AA_LABEL</type>
<position>39.5,-39.5</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>221</ID>
<type>AE_DFF_LOW</type>
<position>30,-448.5</position>
<input>
<ID>IN_0</ID>131 </input>
<output>
<ID>OUTINV_0</ID>130 </output>
<output>
<ID>OUT_0</ID>128 </output>
<input>
<ID>clock</ID>121 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_LABEL</type>
<position>40,-48</position>
<gparam>LABEL_TEXT Q'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>222</ID>
<type>GA_LED</type>
<position>38,-446.5</position>
<input>
<ID>N_in0</ID>128 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>223</ID>
<type>GA_LED</type>
<position>38,-449.5</position>
<input>
<ID>N_in0</ID>130 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>30</ID>
<type>BE_NOR2</type>
<position>8.5,-40</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>10 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>224</ID>
<type>BB_CLOCK</type>
<position>19.5,-452.5</position>
<output>
<ID>CLK</ID>121 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>31</ID>
<type>BE_NOR2</type>
<position>8.5,-48.5</position>
<input>
<ID>IN_0</ID>11 </input>
<input>
<ID>IN_1</ID>9 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>32</ID>
<type>AA_LABEL</type>
<position>0.5,-64</position>
<gparam>LABEL_TEXT SR Flip Flop</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>33</ID>
<type>AA_TOGGLE</type>
<position>-5,-75</position>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>34</ID>
<type>AA_TOGGLE</type>
<position>-5,-86</position>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>228</ID>
<type>AA_TOGGLE</type>
<position>-6,-449</position>
<output>
<ID>OUT_0</ID>129 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>35</ID>
<type>AA_LABEL</type>
<position>-9,-74.5</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>36</ID>
<type>AA_LABEL</type>
<position>-9,-85.5</position>
<gparam>LABEL_TEXT R</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>37</ID>
<type>GA_LED</type>
<position>39.5,-75</position>
<input>
<ID>N_in0</ID>12 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>231</ID>
<type>AA_LABEL</type>
<position>-9.5,-448.5</position>
<gparam>LABEL_TEXT D</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>38</ID>
<type>GA_LED</type>
<position>40,-85</position>
<input>
<ID>N_in0</ID>13 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>232</ID>
<type>AA_LABEL</type>
<position>9.5,-434</position>
<gparam>LABEL_TEXT T to D Flip Flop</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>39</ID>
<type>AA_LABEL</type>
<position>47,-74</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>40</ID>
<type>AA_LABEL</type>
<position>47,-84.5</position>
<gparam>LABEL_TEXT Q'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>234</ID>
<type>AI_XOR2</type>
<position>5.5,-448</position>
<input>
<ID>IN_0</ID>128 </input>
<input>
<ID>IN_1</ID>129 </input>
<output>
<ID>OUT</ID>131 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>42</ID>
<type>BB_CLOCK</type>
<position>-7,-80</position>
<output>
<ID>CLK</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>44</ID>
<type>BA_NAND2</type>
<position>10.5,-75</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>15 </input>
<output>
<ID>OUT</ID>17 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>45</ID>
<type>BA_NAND2</type>
<position>10.5,-85</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>16 </input>
<output>
<ID>OUT</ID>18 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>46</ID>
<type>BA_NAND2</type>
<position>27.5,-75</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>13 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>47</ID>
<type>BA_NAND2</type>
<position>27.5,-85</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>18 </input>
<output>
<ID>OUT</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>48</ID>
<type>AA_LABEL</type>
<position>0,-96</position>
<gparam>LABEL_TEXT D Flip Flop</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>49</ID>
<type>AA_TOGGLE</type>
<position>-7.5,-106.5</position>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>51</ID>
<type>AA_LABEL</type>
<position>-11.5,-106</position>
<gparam>LABEL_TEXT D</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>53</ID>
<type>GA_LED</type>
<position>52,-107.5</position>
<input>
<ID>N_in0</ID>19 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>54</ID>
<type>GA_LED</type>
<position>52.5,-117.5</position>
<input>
<ID>N_in0</ID>20 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>55</ID>
<type>AA_LABEL</type>
<position>59.5,-106.5</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>56</ID>
<type>AA_LABEL</type>
<position>59.5,-117</position>
<gparam>LABEL_TEXT Q'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>57</ID>
<type>BB_CLOCK</type>
<position>5.5,-112.5</position>
<output>
<ID>CLK</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>58</ID>
<type>BA_NAND2</type>
<position>23,-107.5</position>
<input>
<ID>IN_0</ID>21 </input>
<input>
<ID>IN_1</ID>22 </input>
<output>
<ID>OUT</ID>24 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>59</ID>
<type>BA_NAND2</type>
<position>23,-117.5</position>
<input>
<ID>IN_0</ID>22 </input>
<input>
<ID>IN_1</ID>26 </input>
<output>
<ID>OUT</ID>25 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>60</ID>
<type>BA_NAND2</type>
<position>40,-107.5</position>
<input>
<ID>IN_0</ID>24 </input>
<input>
<ID>IN_1</ID>20 </input>
<output>
<ID>OUT</ID>19 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>61</ID>
<type>BA_NAND2</type>
<position>40,-117.5</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>25 </input>
<output>
<ID>OUT</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>63</ID>
<type>AA_INVERTER</type>
<position>-3,-115</position>
<input>
<ID>IN_0</ID>21 </input>
<output>
<ID>OUT_0</ID>26 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>64</ID>
<type>AA_LABEL</type>
<position>5.5,-108</position>
<gparam>LABEL_TEXT Clk</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>65</ID>
<type>AA_LABEL</type>
<position>-13,-79.5</position>
<gparam>LABEL_TEXT Clk</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>66</ID>
<type>AA_LABEL</type>
<position>2,-129.5</position>
<gparam>LABEL_TEXT JK  Flip Flop</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>68</ID>
<type>AE_DFF_LOW</type>
<position>91.5,-111.5</position>
<input>
<ID>IN_0</ID>27 </input>
<output>
<ID>OUTINV_0</ID>30 </output>
<output>
<ID>OUT_0</ID>29 </output>
<input>
<ID>clock</ID>28 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>69</ID>
<type>AA_TOGGLE</type>
<position>83,-109.5</position>
<output>
<ID>OUT_0</ID>27 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>70</ID>
<type>BB_CLOCK</type>
<position>83,-113.5</position>
<output>
<ID>CLK</ID>28 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>71</ID>
<type>GA_LED</type>
<position>98,-109.5</position>
<input>
<ID>N_in0</ID>29 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>72</ID>
<type>GA_LED</type>
<position>98.5,-112.5</position>
<input>
<ID>N_in0</ID>30 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>91</ID>
<type>BE_JKFF_LOW</type>
<position>8.5,-142.5</position>
<input>
<ID>J</ID>42 </input>
<input>
<ID>K</ID>43 </input>
<output>
<ID>Q</ID>45 </output>
<input>
<ID>clock</ID>44 </input>
<output>
<ID>nQ</ID>46 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>93</ID>
<type>AA_TOGGLE</type>
<position>0.5,-140.5</position>
<output>
<ID>OUT_0</ID>42 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>94</ID>
<type>AA_TOGGLE</type>
<position>0.5,-144.5</position>
<output>
<ID>OUT_0</ID>43 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>96</ID>
<type>BB_CLOCK</type>
<position>-6,-142.5</position>
<output>
<ID>CLK</ID>44 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>98</ID>
<type>GA_LED</type>
<position>14.5,-140.5</position>
<input>
<ID>N_in0</ID>45 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>99</ID>
<type>GA_LED</type>
<position>15,-144.5</position>
<input>
<ID>N_in0</ID>46 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>101</ID>
<type>AA_LABEL</type>
<position>21.5,-140</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>102</ID>
<type>AA_LABEL</type>
<position>22,-144</position>
<gparam>LABEL_TEXT Q'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>103</ID>
<type>AA_LABEL</type>
<position>7,-154.5</position>
<gparam>LABEL_TEXT D to SR  Flip Flop</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>105</ID>
<type>AE_DFF_LOW</type>
<position>28,-170.5</position>
<input>
<ID>IN_0</ID>55 </input>
<output>
<ID>OUTINV_0</ID>52 </output>
<output>
<ID>OUT_0</ID>51 </output>
<input>
<ID>clock</ID>47 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>106</ID>
<type>AA_TOGGLE</type>
<position>-10,-165</position>
<output>
<ID>OUT_0</ID>49 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>107</ID>
<type>BB_CLOCK</type>
<position>15.5,-171.5</position>
<output>
<ID>CLK</ID>47 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>108</ID>
<type>AA_TOGGLE</type>
<position>-6.5,-165</position>
<output>
<ID>OUT_0</ID>53 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>110</ID>
<type>AA_INVERTER</type>
<position>-10,-172.5</position>
<input>
<ID>IN_0</ID>49 </input>
<output>
<ID>OUT_0</ID>50 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>112</ID>
<type>AA_AND2</type>
<position>-5,-178</position>
<input>
<ID>IN_0</ID>50 </input>
<input>
<ID>IN_1</ID>51 </input>
<output>
<ID>OUT</ID>54 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>113</ID>
<type>GA_LED</type>
<position>42,-168.5</position>
<input>
<ID>N_in0</ID>51 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>114</ID>
<type>GA_LED</type>
<position>42,-171.5</position>
<input>
<ID>N_in0</ID>52 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>115</ID>
<type>AA_LABEL</type>
<position>46.5,-168</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>116</ID>
<type>AA_LABEL</type>
<position>47,-172</position>
<gparam>LABEL_TEXT Q'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>118</ID>
<type>AE_OR2</type>
<position>4,-168.5</position>
<input>
<ID>IN_0</ID>53 </input>
<input>
<ID>IN_1</ID>54 </input>
<output>
<ID>OUT</ID>55 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>119</ID>
<type>AA_LABEL</type>
<position>-6,-161.5</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>120</ID>
<type>AA_LABEL</type>
<position>-10,-161.5</position>
<gparam>LABEL_TEXT R</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>121</ID>
<type>AA_TOGGLE</type>
<position>-11,-204.5</position>
<output>
<ID>OUT_0</ID>56 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>122</ID>
<type>AA_TOGGLE</type>
<position>-7.5,-204.5</position>
<output>
<ID>OUT_0</ID>58 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>123</ID>
<type>AA_INVERTER</type>
<position>-11,-212</position>
<input>
<ID>IN_0</ID>56 </input>
<output>
<ID>OUT_0</ID>57 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>124</ID>
<type>AA_AND2</type>
<position>-6,-217.5</position>
<input>
<ID>IN_0</ID>57 </input>
<input>
<ID>IN_1</ID>60 </input>
<output>
<ID>OUT</ID>59 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>125</ID>
<type>AE_OR2</type>
<position>3.5,-208</position>
<input>
<ID>IN_0</ID>58 </input>
<input>
<ID>IN_1</ID>59 </input>
<output>
<ID>OUT</ID>65 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>126</ID>
<type>AA_LABEL</type>
<position>-7,-201</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>127</ID>
<type>AA_LABEL</type>
<position>-11,-201</position>
<gparam>LABEL_TEXT R</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>128</ID>
<type>GA_LED</type>
<position>58,-208</position>
<input>
<ID>N_in0</ID>60 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>129</ID>
<type>GA_LED</type>
<position>58.5,-218</position>
<input>
<ID>N_in0</ID>61 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>130</ID>
<type>AA_LABEL</type>
<position>65.5,-207</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>131</ID>
<type>AA_LABEL</type>
<position>65.5,-217.5</position>
<gparam>LABEL_TEXT Q'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>132</ID>
<type>BB_CLOCK</type>
<position>11.5,-213</position>
<output>
<ID>CLK</ID>62 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>133</ID>
<type>BA_NAND2</type>
<position>29,-208</position>
<input>
<ID>IN_0</ID>65 </input>
<input>
<ID>IN_1</ID>62 </input>
<output>
<ID>OUT</ID>63 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>134</ID>
<type>BA_NAND2</type>
<position>29,-222.5</position>
<input>
<ID>IN_0</ID>62 </input>
<input>
<ID>IN_1</ID>66 </input>
<output>
<ID>OUT</ID>64 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>135</ID>
<type>BA_NAND2</type>
<position>46,-208</position>
<input>
<ID>IN_0</ID>63 </input>
<input>
<ID>IN_1</ID>61 </input>
<output>
<ID>OUT</ID>60 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>136</ID>
<type>BA_NAND2</type>
<position>46,-218</position>
<input>
<ID>IN_0</ID>60 </input>
<input>
<ID>IN_1</ID>64 </input>
<output>
<ID>OUT</ID>61 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>137</ID>
<type>AA_LABEL</type>
<position>18,-214.5</position>
<gparam>LABEL_TEXT Clk</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>138</ID>
<type>AA_INVERTER</type>
<position>7.5,-219.5</position>
<input>
<ID>IN_0</ID>65 </input>
<output>
<ID>OUT_0</ID>66 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>139</ID>
<type>AA_LABEL</type>
<position>6.5,-249</position>
<gparam>LABEL_TEXT D to T  Flip Flop</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>140</ID>
<type>AE_DFF_LOW</type>
<position>27.5,-265</position>
<input>
<ID>IN_0</ID>75 </input>
<output>
<ID>OUTINV_0</ID>71 </output>
<output>
<ID>OUT_0</ID>70 </output>
<input>
<ID>clock</ID>67 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>142</ID>
<type>BB_CLOCK</type>
<position>15,-266</position>
<output>
<ID>CLK</ID>67 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>143</ID>
<type>AA_TOGGLE</type>
<position>-7,-259.5</position>
<output>
<ID>OUT_0</ID>77 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>146</ID>
<type>GA_LED</type>
<position>41.5,-263</position>
<input>
<ID>N_in0</ID>70 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>147</ID>
<type>GA_LED</type>
<position>41.5,-266</position>
<input>
<ID>N_in0</ID>71 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>148</ID>
<type>AA_LABEL</type>
<position>46,-262.5</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>149</ID>
<type>AA_LABEL</type>
<position>46.5,-266.5</position>
<gparam>LABEL_TEXT Q'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>151</ID>
<type>AA_LABEL</type>
<position>-7,-255.5</position>
<gparam>LABEL_TEXT T</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>154</ID>
<type>AI_XOR2</type>
<position>4,-263</position>
<input>
<ID>IN_0</ID>70 </input>
<input>
<ID>IN_1</ID>77 </input>
<output>
<ID>OUT</ID>75 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>155</ID>
<type>AA_LABEL</type>
<position>7,-283.5</position>
<gparam>LABEL_TEXT JK to SR  Flip Flop</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>157</ID>
<type>BB_CLOCK</type>
<position>-10,-297.5</position>
<output>
<ID>CLK</ID>86 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>158</ID>
<type>AA_TOGGLE</type>
<position>1.5,-294.5</position>
<output>
<ID>OUT_0</ID>87 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>159</ID>
<type>GA_LED</type>
<position>21.5,-294.5</position>
<input>
<ID>N_in0</ID>84 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>160</ID>
<type>GA_LED</type>
<position>21.5,-298.5</position>
<input>
<ID>N_in0</ID>85 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>161</ID>
<type>AA_LABEL</type>
<position>26,-293.5</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>162</ID>
<type>AA_LABEL</type>
<position>26.5,-298.5</position>
<gparam>LABEL_TEXT Q'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>163</ID>
<type>AA_LABEL</type>
<position>-1.5,-294</position>
<gparam>LABEL_TEXT J</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>166</ID>
<type>BE_JKFF_LOW</type>
<position>11.5,-296.5</position>
<input>
<ID>J</ID>87 </input>
<input>
<ID>K</ID>88 </input>
<output>
<ID>Q</ID>84 </output>
<input>
<ID>clock</ID>86 </input>
<output>
<ID>nQ</ID>85 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>167</ID>
<type>AA_TOGGLE</type>
<position>2,-300.5</position>
<output>
<ID>OUT_0</ID>88 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>168</ID>
<type>AA_LABEL</type>
<position>-1,-300</position>
<gparam>LABEL_TEXT K</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>169</ID>
<type>AA_LABEL</type>
<position>6,-311</position>
<gparam>LABEL_TEXT JK to D  Flip Flop</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>170</ID>
<type>BB_CLOCK</type>
<position>4,-327</position>
<output>
<ID>CLK</ID>91 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>171</ID>
<type>AA_TOGGLE</type>
<position>-9,-320.5</position>
<output>
<ID>OUT_0</ID>94 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>172</ID>
<type>GA_LED</type>
<position>27.5,-327.5</position>
<input>
<ID>N_in0</ID>89 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>173</ID>
<type>GA_LED</type>
<position>27.5,-331.5</position>
<input>
<ID>N_in0</ID>90 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>174</ID>
<type>AA_LABEL</type>
<position>31.5,-327</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>175</ID>
<type>AA_LABEL</type>
<position>32,-331</position>
<gparam>LABEL_TEXT Q'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>176</ID>
<type>AA_LABEL</type>
<position>-9,-317</position>
<gparam>LABEL_TEXT D</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>177</ID>
<type>BE_JKFF_LOW</type>
<position>17.5,-329.5</position>
<input>
<ID>J</ID>94 </input>
<input>
<ID>K</ID>95 </input>
<output>
<ID>Q</ID>89 </output>
<input>
<ID>clock</ID>91 </input>
<output>
<ID>nQ</ID>90 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>181</ID>
<type>AA_INVERTER</type>
<position>-9,-328</position>
<input>
<ID>IN_0</ID>94 </input>
<output>
<ID>OUT_0</ID>95 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>182</ID>
<type>AA_LABEL</type>
<position>7,-341</position>
<gparam>LABEL_TEXT JK to T  Flip Flop</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>183</ID>
<type>BB_CLOCK</type>
<position>4,-353.5</position>
<output>
<ID>CLK</ID>102 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>184</ID>
<type>AA_TOGGLE</type>
<position>-8.5,-355</position>
<output>
<ID>OUT_0</ID>101 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>185</ID>
<type>GA_LED</type>
<position>28.5,-357.5</position>
<input>
<ID>N_in0</ID>96 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>186</ID>
<type>GA_LED</type>
<position>28.5,-361.5</position>
<input>
<ID>N_in0</ID>97 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>187</ID>
<type>AA_LABEL</type>
<position>32.5,-357</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>188</ID>
<type>AA_LABEL</type>
<position>33,-361</position>
<gparam>LABEL_TEXT Q'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>189</ID>
<type>AA_LABEL</type>
<position>-11.5,-354.5</position>
<gparam>LABEL_TEXT T</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>190</ID>
<type>BE_JKFF_LOW</type>
<position>18.5,-359.5</position>
<input>
<ID>J</ID>101 </input>
<input>
<ID>K</ID>101 </input>
<output>
<ID>Q</ID>96 </output>
<input>
<ID>clock</ID>102 </input>
<output>
<ID>nQ</ID>97 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>192</ID>
<type>AA_LABEL</type>
<position>7.5,-372.5</position>
<gparam>LABEL_TEXT T to SR  Flip Flop</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-8.5,-5,-1.5,-5</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<connection>
<GID>10</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-8.5,-15.5,-1.5,-15.5</points>
<connection>
<GID>11</GID>
<name>IN_1</name></connection>
<connection>
<GID>5</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4.5,-6,29.5,-6</points>
<connection>
<GID>10</GID>
<name>OUT</name></connection>
<connection>
<GID>7</GID>
<name>N_in0</name></connection>
<intersection>7 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>7,-13.5,7,-6</points>
<intersection>-13.5 8</intersection>
<intersection>-6 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-1.5,-13.5,7,-13.5</points>
<connection>
<GID>11</GID>
<name>IN_0</name></connection>
<intersection>7 7</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1.5,-14.5,29,-14.5</points>
<connection>
<GID>8</GID>
<name>N_in0</name></connection>
<connection>
<GID>11</GID>
<name>OUT</name></connection>
<intersection>-1.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-1.5,-14.5,-1.5,-7</points>
<connection>
<GID>10</GID>
<name>IN_1</name></connection>
<intersection>-14.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-6,-39,5.5,-39</points>
<connection>
<GID>21</GID>
<name>OUT_0</name></connection>
<connection>
<GID>30</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-6,-49.5,5.5,-49.5</points>
<connection>
<GID>22</GID>
<name>OUT_0</name></connection>
<connection>
<GID>31</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>1,-48.5,31.5,-48.5</points>
<connection>
<GID>31</GID>
<name>OUT</name></connection>
<connection>
<GID>26</GID>
<name>N_in0</name></connection>
<intersection>1 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>1,-48.5,1,-41</points>
<intersection>-48.5 1</intersection>
<intersection>-41 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>1,-41,5.5,-41</points>
<connection>
<GID>30</GID>
<name>IN_1</name></connection>
<intersection>1 4</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>11.5,-40,31.5,-40</points>
<connection>
<GID>25</GID>
<name>N_in0</name></connection>
<connection>
<GID>30</GID>
<name>OUT</name></connection>
<intersection>16 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>16,-47.5,16,-40</points>
<intersection>-47.5 4</intersection>
<intersection>-40 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>5.5,-47.5,16,-47.5</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<intersection>16 3</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-75,38.5,-75</points>
<connection>
<GID>46</GID>
<name>OUT</name></connection>
<connection>
<GID>37</GID>
<name>N_in0</name></connection>
<intersection>32.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>32.5,-84,32.5,-75</points>
<intersection>-84 5</intersection>
<intersection>-75 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>24.5,-84,32.5,-84</points>
<connection>
<GID>47</GID>
<name>IN_0</name></connection>
<intersection>32.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>21.5,-85,39,-85</points>
<connection>
<GID>47</GID>
<name>OUT</name></connection>
<connection>
<GID>38</GID>
<name>N_in0</name></connection>
<intersection>21.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>21.5,-85,21.5,-76</points>
<intersection>-85 1</intersection>
<intersection>-76 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>21.5,-76,24.5,-76</points>
<connection>
<GID>46</GID>
<name>IN_1</name></connection>
<intersection>21.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2,-75,2,-74</points>
<intersection>-75 2</intersection>
<intersection>-74 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>2,-74,7.5,-74</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>2 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-3,-75,2,-75</points>
<connection>
<GID>33</GID>
<name>OUT_0</name></connection>
<intersection>2 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2,-84,2,-76</points>
<intersection>-84 3</intersection>
<intersection>-80 2</intersection>
<intersection>-76 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>2,-76,7.5,-76</points>
<connection>
<GID>44</GID>
<name>IN_1</name></connection>
<intersection>2 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-3,-80,2,-80</points>
<connection>
<GID>42</GID>
<name>CLK</name></connection>
<intersection>2 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>2,-84,7.5,-84</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<intersection>2 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-3,-86,7.5,-86</points>
<connection>
<GID>45</GID>
<name>IN_1</name></connection>
<connection>
<GID>34</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19,-75,19,-74</points>
<intersection>-75 2</intersection>
<intersection>-74 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>19,-74,24.5,-74</points>
<connection>
<GID>46</GID>
<name>IN_0</name></connection>
<intersection>19 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13.5,-75,19,-75</points>
<connection>
<GID>44</GID>
<name>OUT</name></connection>
<intersection>19 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19,-86,19,-85</points>
<intersection>-86 1</intersection>
<intersection>-85 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>19,-86,24.5,-86</points>
<connection>
<GID>47</GID>
<name>IN_1</name></connection>
<intersection>19 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13.5,-85,19,-85</points>
<connection>
<GID>45</GID>
<name>OUT</name></connection>
<intersection>19 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>43,-107.5,51,-107.5</points>
<connection>
<GID>53</GID>
<name>N_in0</name></connection>
<connection>
<GID>60</GID>
<name>OUT</name></connection>
<intersection>45.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>45.5,-116.5,45.5,-107.5</points>
<intersection>-116.5 5</intersection>
<intersection>-107.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>37,-116.5,45.5,-116.5</points>
<connection>
<GID>61</GID>
<name>IN_0</name></connection>
<intersection>45.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,-117.5,51.5,-117.5</points>
<connection>
<GID>54</GID>
<name>N_in0</name></connection>
<connection>
<GID>61</GID>
<name>OUT</name></connection>
<intersection>34 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>34,-117.5,34,-108.5</points>
<intersection>-117.5 1</intersection>
<intersection>-108.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>34,-108.5,37,-108.5</points>
<connection>
<GID>60</GID>
<name>IN_1</name></connection>
<intersection>34 6</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-5.5,-106.5,20,-106.5</points>
<connection>
<GID>49</GID>
<name>OUT_0</name></connection>
<connection>
<GID>58</GID>
<name>IN_0</name></connection>
<intersection>-3 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-3,-112,-3,-106.5</points>
<connection>
<GID>63</GID>
<name>IN_0</name></connection>
<intersection>-106.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14.5,-116.5,14.5,-108.5</points>
<intersection>-116.5 3</intersection>
<intersection>-112.5 2</intersection>
<intersection>-108.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>14.5,-108.5,20,-108.5</points>
<connection>
<GID>58</GID>
<name>IN_1</name></connection>
<intersection>14.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>9.5,-112.5,14.5,-112.5</points>
<connection>
<GID>57</GID>
<name>CLK</name></connection>
<intersection>14.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>14.5,-116.5,20,-116.5</points>
<connection>
<GID>59</GID>
<name>IN_0</name></connection>
<intersection>14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,-107.5,31.5,-106.5</points>
<intersection>-107.5 2</intersection>
<intersection>-106.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31.5,-106.5,37,-106.5</points>
<connection>
<GID>60</GID>
<name>IN_0</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-107.5,31.5,-107.5</points>
<connection>
<GID>58</GID>
<name>OUT</name></connection>
<intersection>31.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,-118.5,31.5,-117.5</points>
<intersection>-118.5 1</intersection>
<intersection>-117.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31.5,-118.5,37,-118.5</points>
<connection>
<GID>61</GID>
<name>IN_1</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-117.5,31.5,-117.5</points>
<connection>
<GID>59</GID>
<name>OUT</name></connection>
<intersection>31.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-3,-118.5,20,-118.5</points>
<connection>
<GID>59</GID>
<name>IN_1</name></connection>
<intersection>-3 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-3,-118.5,-3,-118</points>
<connection>
<GID>63</GID>
<name>OUT_0</name></connection>
<intersection>-118.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>85,-109.5,88.5,-109.5</points>
<connection>
<GID>68</GID>
<name>IN_0</name></connection>
<connection>
<GID>69</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87.5,-113.5,87.5,-112.5</points>
<intersection>-113.5 2</intersection>
<intersection>-112.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>87.5,-112.5,88.5,-112.5</points>
<connection>
<GID>68</GID>
<name>clock</name></connection>
<intersection>87.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>87,-113.5,87.5,-113.5</points>
<connection>
<GID>70</GID>
<name>CLK</name></connection>
<intersection>87.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>94.5,-109.5,97,-109.5</points>
<connection>
<GID>71</GID>
<name>N_in0</name></connection>
<connection>
<GID>68</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>94.5,-112.5,97.5,-112.5</points>
<connection>
<GID>72</GID>
<name>N_in0</name></connection>
<connection>
<GID>68</GID>
<name>OUTINV_0</name></connection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>2.5,-140.5,5.5,-140.5</points>
<connection>
<GID>91</GID>
<name>J</name></connection>
<connection>
<GID>93</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>2.5,-144.5,5.5,-144.5</points>
<connection>
<GID>94</GID>
<name>OUT_0</name></connection>
<intersection>5.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>5.5,-144.5,5.5,-144.5</points>
<connection>
<GID>91</GID>
<name>K</name></connection>
<intersection>-144.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-2,-142.5,5.5,-142.5</points>
<connection>
<GID>91</GID>
<name>clock</name></connection>
<connection>
<GID>96</GID>
<name>CLK</name></connection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>11.5,-140.5,13.5,-140.5</points>
<connection>
<GID>98</GID>
<name>N_in0</name></connection>
<connection>
<GID>91</GID>
<name>Q</name></connection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>11.5,-144.5,14,-144.5</points>
<connection>
<GID>99</GID>
<name>N_in0</name></connection>
<connection>
<GID>91</GID>
<name>nQ</name></connection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-171.5,25,-171.5</points>
<connection>
<GID>105</GID>
<name>clock</name></connection>
<connection>
<GID>107</GID>
<name>CLK</name></connection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-10,-169.5,-10,-167</points>
<connection>
<GID>106</GID>
<name>OUT_0</name></connection>
<connection>
<GID>110</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-10,-177,-10,-175.5</points>
<connection>
<GID>110</GID>
<name>OUT_0</name></connection>
<intersection>-177 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-10,-177,-8,-177</points>
<connection>
<GID>112</GID>
<name>IN_0</name></connection>
<intersection>-10 0</intersection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-8,-179,39,-179</points>
<connection>
<GID>112</GID>
<name>IN_1</name></connection>
<intersection>39 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>39,-179,39,-168.5</points>
<intersection>-179 1</intersection>
<intersection>-168.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>31,-168.5,41,-168.5</points>
<connection>
<GID>105</GID>
<name>OUT_0</name></connection>
<connection>
<GID>113</GID>
<name>N_in0</name></connection>
<intersection>39 4</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31,-171.5,41,-171.5</points>
<connection>
<GID>105</GID>
<name>OUTINV_0</name></connection>
<connection>
<GID>114</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-6.5,-167.5,-6.5,-167</points>
<connection>
<GID>108</GID>
<name>OUT_0</name></connection>
<intersection>-167.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-6.5,-167.5,1,-167.5</points>
<connection>
<GID>118</GID>
<name>IN_0</name></connection>
<intersection>-6.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-0.5,-178,-0.5,-169.5</points>
<intersection>-178 2</intersection>
<intersection>-169.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-0.5,-169.5,1,-169.5</points>
<connection>
<GID>118</GID>
<name>IN_1</name></connection>
<intersection>-0.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-2,-178,-0.5,-178</points>
<connection>
<GID>112</GID>
<name>OUT</name></connection>
<intersection>-0.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7,-168.5,25,-168.5</points>
<connection>
<GID>105</GID>
<name>IN_0</name></connection>
<connection>
<GID>118</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-11,-209,-11,-206.5</points>
<connection>
<GID>123</GID>
<name>IN_0</name></connection>
<connection>
<GID>121</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-11,-216.5,-11,-215</points>
<connection>
<GID>123</GID>
<name>OUT_0</name></connection>
<intersection>-216.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-11,-216.5,-9,-216.5</points>
<connection>
<GID>124</GID>
<name>IN_0</name></connection>
<intersection>-11 0</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-7.5,-207,-7.5,-206.5</points>
<connection>
<GID>122</GID>
<name>OUT_0</name></connection>
<intersection>-207 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-7.5,-207,0.5,-207</points>
<connection>
<GID>125</GID>
<name>IN_0</name></connection>
<intersection>-7.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1.5,-217.5,-1.5,-209</points>
<intersection>-217.5 2</intersection>
<intersection>-209 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1.5,-209,0.5,-209</points>
<connection>
<GID>125</GID>
<name>IN_1</name></connection>
<intersection>-1.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-3,-217.5,-1.5,-217.5</points>
<connection>
<GID>124</GID>
<name>OUT</name></connection>
<intersection>-1.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>49,-208,57,-208</points>
<connection>
<GID>135</GID>
<name>OUT</name></connection>
<connection>
<GID>128</GID>
<name>N_in0</name></connection>
<intersection>51.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>51.5,-231,51.5,-208</points>
<intersection>-231 5</intersection>
<intersection>-208 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-9,-231,51.5,-231</points>
<intersection>-9 8</intersection>
<intersection>43 9</intersection>
<intersection>51.5 4</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-9,-231,-9,-218.5</points>
<connection>
<GID>124</GID>
<name>IN_1</name></connection>
<intersection>-231 5</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>43,-231,43,-217</points>
<connection>
<GID>136</GID>
<name>IN_0</name></connection>
<intersection>-231 5</intersection></vsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40,-218,57.5,-218</points>
<connection>
<GID>136</GID>
<name>OUT</name></connection>
<connection>
<GID>129</GID>
<name>N_in0</name></connection>
<intersection>40 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>40,-218,40,-209</points>
<intersection>-218 1</intersection>
<intersection>-209 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>40,-209,43,-209</points>
<connection>
<GID>135</GID>
<name>IN_1</name></connection>
<intersection>40 6</intersection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,-221.5,20.5,-209</points>
<intersection>-221.5 3</intersection>
<intersection>-213 2</intersection>
<intersection>-209 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20.5,-209,26,-209</points>
<connection>
<GID>133</GID>
<name>IN_1</name></connection>
<intersection>20.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>15.5,-213,20.5,-213</points>
<connection>
<GID>132</GID>
<name>CLK</name></connection>
<intersection>20.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>20.5,-221.5,26,-221.5</points>
<connection>
<GID>134</GID>
<name>IN_0</name></connection>
<intersection>20.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37.5,-208,37.5,-207</points>
<intersection>-208 2</intersection>
<intersection>-207 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37.5,-207,43,-207</points>
<connection>
<GID>135</GID>
<name>IN_0</name></connection>
<intersection>37.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32,-208,37.5,-208</points>
<connection>
<GID>133</GID>
<name>OUT</name></connection>
<intersection>37.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37.5,-222.5,37.5,-219</points>
<intersection>-222.5 2</intersection>
<intersection>-219 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37.5,-219,43,-219</points>
<connection>
<GID>136</GID>
<name>IN_1</name></connection>
<intersection>37.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32,-222.5,37.5,-222.5</points>
<connection>
<GID>134</GID>
<name>OUT</name></connection>
<intersection>37.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16,-208,16,-207</points>
<intersection>-208 2</intersection>
<intersection>-207 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>16,-207,26,-207</points>
<connection>
<GID>133</GID>
<name>IN_0</name></connection>
<intersection>16 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>6.5,-208,16,-208</points>
<connection>
<GID>125</GID>
<name>OUT</name></connection>
<intersection>7.5 3</intersection>
<intersection>16 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>7.5,-216.5,7.5,-208</points>
<connection>
<GID>138</GID>
<name>IN_0</name></connection>
<intersection>-208 2</intersection></vsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7.5,-223.5,7.5,-222.5</points>
<connection>
<GID>138</GID>
<name>OUT_0</name></connection>
<intersection>-223.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>7.5,-223.5,26,-223.5</points>
<connection>
<GID>134</GID>
<name>IN_1</name></connection>
<intersection>7.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19,-266,24.5,-266</points>
<connection>
<GID>142</GID>
<name>CLK</name></connection>
<connection>
<GID>140</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<hsegment>
<ID>9</ID>
<points>1,-258,40.5,-258</points>
<intersection>1 10</intersection>
<intersection>30.5 14</intersection>
<intersection>40.5 12</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>1,-262,1,-258</points>
<connection>
<GID>154</GID>
<name>IN_0</name></connection>
<intersection>-258 9</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>40.5,-263,40.5,-258</points>
<connection>
<GID>146</GID>
<name>N_in0</name></connection>
<intersection>-258 9</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>30.5,-263,30.5,-258</points>
<connection>
<GID>140</GID>
<name>OUT_0</name></connection>
<intersection>-258 9</intersection></vsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-266,40.5,-266</points>
<connection>
<GID>147</GID>
<name>N_in0</name></connection>
<connection>
<GID>140</GID>
<name>OUTINV_0</name></connection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7,-263,24.5,-263</points>
<connection>
<GID>140</GID>
<name>IN_0</name></connection>
<connection>
<GID>154</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-7,-264,-7,-261.5</points>
<connection>
<GID>143</GID>
<name>OUT_0</name></connection>
<intersection>-264 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-7,-264,1,-264</points>
<connection>
<GID>154</GID>
<name>IN_1</name></connection>
<intersection>-7 0</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>14.5,-294.5,20.5,-294.5</points>
<connection>
<GID>159</GID>
<name>N_in0</name></connection>
<connection>
<GID>166</GID>
<name>Q</name></connection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>14.5,-298.5,20.5,-298.5</points>
<connection>
<GID>160</GID>
<name>N_in0</name></connection>
<connection>
<GID>166</GID>
<name>nQ</name></connection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3.5,-297.5,3.5,-296.5</points>
<intersection>-297.5 2</intersection>
<intersection>-296.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>3.5,-296.5,8.5,-296.5</points>
<connection>
<GID>166</GID>
<name>clock</name></connection>
<intersection>3.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-6,-297.5,3.5,-297.5</points>
<connection>
<GID>157</GID>
<name>CLK</name></connection>
<intersection>3.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3.5,-294.5,8.5,-294.5</points>
<connection>
<GID>158</GID>
<name>OUT_0</name></connection>
<connection>
<GID>166</GID>
<name>J</name></connection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6,-300.5,6,-298.5</points>
<intersection>-300.5 2</intersection>
<intersection>-298.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>6,-298.5,8.5,-298.5</points>
<connection>
<GID>166</GID>
<name>K</name></connection>
<intersection>6 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>4,-300.5,6,-300.5</points>
<connection>
<GID>167</GID>
<name>OUT_0</name></connection>
<intersection>6 0</intersection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<hsegment>
<ID>14</ID>
<points>20.5,-327.5,26.5,-327.5</points>
<connection>
<GID>172</GID>
<name>N_in0</name></connection>
<connection>
<GID>177</GID>
<name>Q</name></connection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<hsegment>
<ID>14</ID>
<points>20.5,-331.5,26.5,-331.5</points>
<connection>
<GID>173</GID>
<name>N_in0</name></connection>
<connection>
<GID>177</GID>
<name>nQ</name></connection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>8,-329.5,14.5,-329.5</points>
<connection>
<GID>177</GID>
<name>clock</name></connection>
<intersection>8 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>8,-329.5,8,-327</points>
<connection>
<GID>170</GID>
<name>CLK</name></connection>
<intersection>-329.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-9,-325,-9,-322.5</points>
<connection>
<GID>171</GID>
<name>OUT_0</name></connection>
<connection>
<GID>181</GID>
<name>IN_0</name></connection>
<intersection>-324 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-9,-324,14.5,-324</points>
<intersection>-9 0</intersection>
<intersection>14.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>14.5,-327.5,14.5,-324</points>
<connection>
<GID>177</GID>
<name>J</name></connection>
<intersection>-324 3</intersection></vsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-9,-331.5,-9,-331</points>
<connection>
<GID>181</GID>
<name>OUT_0</name></connection>
<intersection>-331.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-9,-331.5,14.5,-331.5</points>
<connection>
<GID>177</GID>
<name>K</name></connection>
<intersection>-9 0</intersection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<hsegment>
<ID>14</ID>
<points>21.5,-357.5,27.5,-357.5</points>
<connection>
<GID>185</GID>
<name>N_in0</name></connection>
<connection>
<GID>190</GID>
<name>Q</name></connection></hsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<hsegment>
<ID>14</ID>
<points>21.5,-361.5,27.5,-361.5</points>
<connection>
<GID>186</GID>
<name>N_in0</name></connection>
<connection>
<GID>190</GID>
<name>nQ</name></connection></hsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-6.5,-355,-3.5,-355</points>
<connection>
<GID>184</GID>
<name>OUT_0</name></connection>
<intersection>-3.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-3.5,-361.5,-3.5,-355</points>
<intersection>-361.5 6</intersection>
<intersection>-357.5 7</intersection>
<intersection>-355 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-3.5,-361.5,15.5,-361.5</points>
<connection>
<GID>190</GID>
<name>K</name></connection>
<intersection>-3.5 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-3.5,-357.5,15.5,-357.5</points>
<connection>
<GID>190</GID>
<name>J</name></connection>
<intersection>-3.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11.5,-359.5,11.5,-353.5</points>
<intersection>-359.5 2</intersection>
<intersection>-353.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8,-353.5,11.5,-353.5</points>
<connection>
<GID>183</GID>
<name>CLK</name></connection>
<intersection>11.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11.5,-359.5,15.5,-359.5</points>
<connection>
<GID>190</GID>
<name>clock</name></connection>
<intersection>11.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1.5,-381,35,-381</points>
<intersection>-1.5 3</intersection>
<intersection>31 5</intersection>
<intersection>35 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-1.5,-383,-1.5,-381</points>
<connection>
<GID>200</GID>
<name>IN_0</name></connection>
<intersection>-381 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>35,-385,35,-381</points>
<connection>
<GID>196</GID>
<name>N_in0</name></connection>
<intersection>-381 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>31,-385,31,-381</points>
<connection>
<GID>194</GID>
<name>OUT_0</name></connection>
<intersection>-381 1</intersection></vsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1.5,-397.5,35,-397.5</points>
<intersection>-1.5 4</intersection>
<intersection>31 5</intersection>
<intersection>35 6</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-1.5,-397.5,-1.5,-392.5</points>
<connection>
<GID>201</GID>
<name>IN_1</name></connection>
<intersection>-397.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>31,-397.5,31,-388</points>
<connection>
<GID>194</GID>
<name>OUTINV_0</name></connection>
<intersection>-397.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>35,-397.5,35,-388</points>
<connection>
<GID>197</GID>
<name>N_in0</name></connection>
<intersection>-397.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>21.5,-391,25,-391</points>
<connection>
<GID>198</GID>
<name>CLK</name></connection>
<intersection>25 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>25,-391,25,-388</points>
<connection>
<GID>194</GID>
<name>clock</name></connection>
<intersection>-391 1</intersection></vsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6,-386,6,-384</points>
<intersection>-386 1</intersection>
<intersection>-384 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>6,-386,7,-386</points>
<connection>
<GID>203</GID>
<name>IN_0</name></connection>
<intersection>6 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>4.5,-384,6,-384</points>
<connection>
<GID>200</GID>
<name>OUT</name></connection>
<intersection>6 0</intersection></hsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6,-391.5,6,-388</points>
<intersection>-391.5 2</intersection>
<intersection>-388 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>6,-388,7,-388</points>
<connection>
<GID>203</GID>
<name>IN_1</name></connection>
<intersection>6 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>4.5,-391.5,6,-391.5</points>
<connection>
<GID>201</GID>
<name>OUT</name></connection>
<intersection>6 0</intersection></hsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19,-387,19,-385</points>
<intersection>-387 2</intersection>
<intersection>-385 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>19,-385,25,-385</points>
<connection>
<GID>194</GID>
<name>IN_0</name></connection>
<intersection>19 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13,-387,19,-387</points>
<connection>
<GID>203</GID>
<name>OUT</name></connection>
<intersection>19 0</intersection></hsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-5.5,-385,-1.5,-385</points>
<connection>
<GID>200</GID>
<name>IN_1</name></connection>
<connection>
<GID>205</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-5.5,-390.5,-1.5,-390.5</points>
<connection>
<GID>201</GID>
<name>IN_0</name></connection>
<connection>
<GID>206</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1.5,-409.5,35,-409.5</points>
<intersection>-1.5 3</intersection>
<intersection>31 5</intersection>
<intersection>35 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-1.5,-411.5,-1.5,-409.5</points>
<connection>
<GID>213</GID>
<name>IN_0</name></connection>
<intersection>-409.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>35,-413.5,35,-409.5</points>
<connection>
<GID>210</GID>
<name>N_in0</name></connection>
<intersection>-409.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>31,-413.5,31,-409.5</points>
<connection>
<GID>209</GID>
<name>OUT_0</name></connection>
<intersection>-409.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1.5,-426,35,-426</points>
<intersection>-1.5 4</intersection>
<intersection>31 5</intersection>
<intersection>35 6</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-1.5,-426,-1.5,-421</points>
<connection>
<GID>214</GID>
<name>IN_1</name></connection>
<intersection>-426 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>31,-426,31,-416.5</points>
<connection>
<GID>209</GID>
<name>OUTINV_0</name></connection>
<intersection>-426 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>35,-426,35,-416.5</points>
<connection>
<GID>211</GID>
<name>N_in0</name></connection>
<intersection>-426 1</intersection></vsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>21.5,-419.5,25,-419.5</points>
<connection>
<GID>212</GID>
<name>CLK</name></connection>
<intersection>25 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>25,-419.5,25,-416.5</points>
<connection>
<GID>209</GID>
<name>clock</name></connection>
<intersection>-419.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6,-414.5,6,-412.5</points>
<intersection>-414.5 1</intersection>
<intersection>-412.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>6,-414.5,7,-414.5</points>
<connection>
<GID>215</GID>
<name>IN_0</name></connection>
<intersection>6 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>4.5,-412.5,6,-412.5</points>
<connection>
<GID>213</GID>
<name>OUT</name></connection>
<intersection>6 0</intersection></hsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6,-420,6,-416.5</points>
<intersection>-420 2</intersection>
<intersection>-416.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>6,-416.5,7,-416.5</points>
<connection>
<GID>215</GID>
<name>IN_1</name></connection>
<intersection>6 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>4.5,-420,6,-420</points>
<connection>
<GID>214</GID>
<name>OUT</name></connection>
<intersection>6 0</intersection></hsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19,-415.5,19,-413.5</points>
<intersection>-415.5 2</intersection>
<intersection>-413.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>19,-413.5,25,-413.5</points>
<connection>
<GID>209</GID>
<name>IN_0</name></connection>
<intersection>19 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13,-415.5,19,-415.5</points>
<connection>
<GID>215</GID>
<name>OUT</name></connection>
<intersection>19 0</intersection></hsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-5.5,-413.5,-1.5,-413.5</points>
<connection>
<GID>216</GID>
<name>OUT_0</name></connection>
<connection>
<GID>213</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-5.5,-419,-1.5,-419</points>
<connection>
<GID>217</GID>
<name>OUT_0</name></connection>
<connection>
<GID>214</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>23.5,-452.5,27,-452.5</points>
<connection>
<GID>224</GID>
<name>CLK</name></connection>
<intersection>27 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>27,-452.5,27,-449.5</points>
<connection>
<GID>221</GID>
<name>clock</name></connection>
<intersection>-452.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>2.5,-443.5,37,-443.5</points>
<intersection>2.5 3</intersection>
<intersection>33 5</intersection>
<intersection>37 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>2.5,-447,2.5,-443.5</points>
<connection>
<GID>234</GID>
<name>IN_0</name></connection>
<intersection>-443.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>37,-446.5,37,-443.5</points>
<connection>
<GID>222</GID>
<name>N_in0</name></connection>
<intersection>-443.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>33,-446.5,33,-443.5</points>
<connection>
<GID>221</GID>
<name>OUT_0</name></connection>
<intersection>-443.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-4,-449,2.5,-449</points>
<connection>
<GID>234</GID>
<name>IN_1</name></connection>
<connection>
<GID>228</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>33,-449.5,37,-449.5</points>
<connection>
<GID>223</GID>
<name>N_in0</name></connection>
<connection>
<GID>221</GID>
<name>OUTINV_0</name></connection></hsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17.5,-448,17.5,-446.5</points>
<intersection>-448 2</intersection>
<intersection>-446.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17.5,-446.5,27,-446.5</points>
<connection>
<GID>221</GID>
<name>IN_0</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8.5,-448,17.5,-448</points>
<connection>
<GID>234</GID>
<name>OUT</name></connection>
<intersection>17.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 1>
<page 2>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 2>
<page 3>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 3>
<page 4>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 4>
<page 5>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 5>
<page 6>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 6>
<page 7>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 7>
<page 8>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 8>
<page 9>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 9></circuit>